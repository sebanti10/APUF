`ifndef parameters
`define parameters

    parameter C_LENGTH = 3; //the length of the chain of multiplexer
    
`endif